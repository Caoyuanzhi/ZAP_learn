`include "my_if.sv"
`include "my_transcation.sv"
`include "my_driver.sv"
`include "my_monitor.sv"
//add a confilct on branch
`include "my_env.sv"
`include "assertion/ast_test.sv"
